`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/23/2021 01:46:20 PM
// Design Name: 
// Module Name: PE
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "global.v"

module PE #(
    parameter   KERNEL_SIZE = `KERNEL_SIZE,
    parameter   FM_SIZE     = `FM_SIZE,
    parameter   PADDING     = `PADDING,
    parameter   STRIDE      = `STRIDE,
    localparam  OUT_SIZE    = ((FM_SIZE - KERNEL_SIZE + 2 * PADDING) / STRIDE) + 1
)(
    input wire i_clk,
    input wire i_en,
    input wire signed [`A_DSP_WIDTH-1:0]        i_data,
    input wire signed [`B_DSP_WIDTH-1:0]        i_weight,
    input wire signed [`OUTPUT_DSP_WIDTH-1:0]   i_partoutvalue,

    output wire o_en,
    output wire signed [`OUTPUT_DSP_WIDTH-1:0] o_data
);
    assign o_en = i_en;


    DSP48E1 #(
        // Feature Control Attributes: Data Path Selection
        .A_INPUT("DIRECT"),                 // Selects A input source, "DIRECT" (A port) or "CASCADE" (ACIN port)
        .B_INPUT("DIRECT"),                 // Selects B input source, "DIRECT" (B port) or "CASCADE" (BCIN port)
        .USE_DPORT("FALSE"),                // Select D port usage (TRUE or FALSE)
        .USE_MULT("MULTIPLY"),              // Select multiplier usage ("MULTIPLY", "DYNAMIC", or "NONE")
        .USE_SIMD("ONE48"),                 // SIMD selection ("ONE48", "TWO24", "FOUR12")

        // Pattern Detector Attributes: Pattern Detection Configuration
        .AUTORESET_PATDET("NO_RESET"),      // "NO_RESET", "RESET_MATCH", "RESET_NOT_MATCH" 
        .MASK(48'h3fffffffffff),            // 48-bit mask value for pattern detect (1=ignore)
        .PATTERN(48'h000000000000),         // 48-bit pattern match for pattern detect
        .SEL_MASK("MASK"),                  // "C", "MASK", "ROUNDING_MODE1", "ROUNDING_MODE2" 
        .SEL_PATTERN("PATTERN"),            // Select pattern value ("PATTERN" or "C")
        .USE_PATTERN_DETECT("NO_PATDET"),   // Enable pattern detect ("PATDET" or "NO_PATDET")

        // Register Control Attributes: Pipeline Register Configuration
        .ACASCREG(0),                       // Number of pipeline stages between A/ACIN and ACOUT (0, 1 or 2)
        .ADREG(0),                          // Number of pipeline stages for pre-adder (0 or 1)
        .ALUMODEREG(0),                     // Number of pipeline stages for ALUMODE (0 or 1)
        .AREG(0),                           // Number of pipeline stages for A (0, 1 or 2)
        .BCASCREG(0),                       // Number of pipeline stages between B/BCIN and BCOUT (0, 1 or 2)
        .BREG(0),                           // Number of pipeline stages for B (0, 1 or 2)
        .CARRYINREG(0),                     // Number of pipeline stages for CARRYIN (0 or 1)
        .CARRYINSELREG(0),                  // Number of pipeline stages for CARRYINSEL (0 or 1)
        .CREG(0),                           // Number of pipeline stages for C (0 or 1)
        .DREG(0),                           // Number of pipeline stages for D (0 or 1)
        .INMODEREG(0),                      // Number of pipeline stages for INMODE (0 or 1)
        .MREG(0),                           // Number of multiplier pipeline stages (0 or 1)
        .OPMODEREG(0),                      // Number of pipeline stages for OPMODE (0 or 1)
        .PREG(0)                            // Number of pipeline stages for P (0 or 1)
    )
    DSP48E1_inst (
        // Cascade: 30-bit (each) output: Cascade Ports
        .ACOUT(),                           // 30-bit output: A port cascade output
        .BCOUT(),                           // 18-bit output: B port cascade output
        .CARRYCASCOUT(),                    // 1-bit output: Cascade carry output
        .MULTSIGNOUT(),                     // 1-bit output: Multiplier sign cascade output
        .PCOUT(),                           // 48-bit output: Cascade output

        // Control: 1-bit (each) output: Control Inputs/Status Bits
        .OVERFLOW(),                        // 1-bit output: Overflow in add/acc output
        .PATTERNBDETECT(),                  // 1-bit output: Pattern bar detect output
        .PATTERNDETECT(),                   // 1-bit output: Pattern detect output
        .UNDERFLOW(),                       // 1-bit output: Underflow in add/acc output

        // Data: 4-bit (each) output: Data Ports
        .CARRYOUT(),                        // 4-bit output: Carry output
        .P(o_data),                         // 48-bit output: Primary data output

        // Cascade: 30-bit (each) input: Cascade Ports
        .ACIN(0),                           // 30-bit input: A cascade data input
        .BCIN(0),                           // 18-bit input: B cascade input
        .CARRYCASCIN(0),                    // 1-bit input: Cascade carry input
        .MULTSIGNIN(0),                     // 1-bit input: Multiplier sign input
        .PCIN(0),                           // 48-bit input: P cascade input

        // Control: 4-bit (each) input: Control Inputs/Status Bits
        .ALUMODE(4'd0),                     // 4-bit input: ALU control input
        .CARRYINSEL(3'd0),                  // 3-bit input: Carry select input
        .CLK(i_clk),                        // 1-bit input: Clock input
        .INMODE(5'd0),                      // 5-bit input: INMODE control input
        .OPMODE(9'b000110101),              // 7-bit input: Operation mode input

        // Data: 30-bit (each) input: Data Ports
        .A(i_data),                         // 30-bit input: A data input
        .B(i_weight),                       // 18-bit input: B data input
        .C(i_partoutvalue),                 // 48-bit input: C data input
        .CARRYIN(0),                        // 1-bit input: Carry input signal
        .D(0),                              // 25-bit input: D data input

        // Reset/Clock Enable: 1-bit (each) input: Reset/Clock Enable Inputs
        .CEA1(1),                           // 1-bit input: Clock enable input for 1st stage AREG
        .CEA2(1),                           // 1-bit input: Clock enable input for 2nd stage AREG
        .CEAD(1),                           // 1-bit input: Clock enable input for ADREG
        .CEALUMODE(1),                      // 1-bit input: Clock enable input for ALUMODE
        .CEB1(1),                           // 1-bit input: Clock enable input for 1st stage BREG
        .CEB2(1),                           // 1-bit input: Clock enable input for 2nd stage BREG
        .CEC(1),                            // 1-bit input: Clock enable input for CREG
        .CECARRYIN(1),                      // 1-bit input: Clock enable input for CARRYINREG
        .CECTRL(1),                         // 1-bit input: Clock enable input for OPMODEREG and CARRYINSELREG
        .CED(1),                            // 1-bit input: Clock enable input for DREG
        .CEINMODE(1),                       // 1-bit input: Clock enable input for INMODEREG
        .CEM(1),                            // 1-bit input: Clock enable input for MREG
        .CEP(1),                            // 1-bit input: Clock enable input for PREG
        .RSTA(0),                           // 1-bit input: Reset input for AREG
        .RSTALLCARRYIN(0),                  // 1-bit input: Reset input for CARRYINREG
        .RSTALUMODE(0),                     // 1-bit input: Reset input for ALUMODEREG
        .RSTB(0),                           // 1-bit input: Reset input for BREG
        .RSTC(0),                           // 1-bit input: Reset input for CREG
        .RSTCTRL(0),                        // 1-bit input: Reset input for OPMODEREG and CARRYINSELREG
        .RSTD(0),                           // 1-bit input: Reset input for DREG and ADREG
        .RSTINMODE(0),                      // 1-bit input: Reset input for INMODEREG
        .RSTM(0),                           // 1-bit input: Reset input for MREG
        .RSTP(0)                            // 1-bit input: Reset input for PREG
    );
endmodule
